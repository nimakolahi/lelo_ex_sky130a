*cicsimgen tran

.param SEED=0

*Nothing here

.param mc_mm_switch=0
.param mc_pr_switch=0
.include "/opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_01v8__tt.pm3.spice"
.include "/opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_01v8__mismatch.corner.spice"
.include "/opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8__tt.corner.spice"
.include "/opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8__mismatch.corner.spice"
.include "/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/corners/tt/nonfet.spice"
.include "/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/all.spice"
.include "/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice"
.include "/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice"
.include "/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice"

.lib "../../../tech/ngspice/temperature.spi" Tt

.lib "../../../tech/ngspice/supply.spi" Vt

*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../../work/xsch/LELO_EX.spice
 
*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
IBP 0 IBPS_5U dc 5u
V0  IBNS_20U 0 dc 1
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
*XDUT IBPS_5U VSS IBNS_20U  LELO_EX


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
*.save all
.save i(V0) v(IBPS_5U)


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


tran 1n 10n 1p
write
quit


.endc

.end

