* NGSPICE file created from LELO_EX.ext - technology: sky130A

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt LELO_EX IBPS_5U VSS IBNS_20U
*.subckt LELO_EX IBPS_5U IBNS_20U VSS
X0 IBNS_20U IBPS_5U VSS VSS sky130_fd_pr__nfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X1 IBPS_5U IBPS_5U VSS VSS sky130_fd_pr__nfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X2 VSS IBPS_5U IBNS_20U VSS sky130_fd_pr__nfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X3 IBNS_20U IBPS_5U VSS VSS sky130_fd_pr__nfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X4 IBNS_20U IBPS_5U VSS VSS sky130_fd_pr__nfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X5 VSS IBPS_5U IBNS_20U VSS sky130_fd_pr__nfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X6 VSS IBPS_5U IBPS_5U VSS sky130_fd_pr__nfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X7 VSS IBPS_5U IBNS_20U VSS sky130_fd_pr__nfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X8 IBNS_20U IBPS_5U VSS VSS sky130_fd_pr__nfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X9 VSS IBPS_5U IBNS_20U VSS sky130_fd_pr__nfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
C0 a_n440_286# IBPS_5U 0.15824f
C1 a_n440_n514# IBPS_5U 0.14444f
C2 a_n441_1887# IBPS_5U 0.14406f
C3 IBPS_5U a_n440_n1313# 0.07043f
C4 IBNS_20U a_n440_286# 0.02796f
C5 IBPS_5U a_n441_2690# 0.07043f
C6 a_n441_1087# IBPS_5U 0.16112f
C7 IBNS_20U a_n440_n514# 0.04156f
C8 IBNS_20U a_n441_1887# 0.04251f
C9 IBNS_20U a_n440_n1313# 0.01909f
C10 IBNS_20U a_n441_1087# 0.02169f
C11 IBNS_20U a_n441_2690# 0.02152f
C12 IBNS_20U IBPS_5U 2.30691f
C13 IBNS_20U VSS 4.53066f
C14 IBPS_5U VSS 13.7027f
C15 a_n440_n1313# VSS 0.67275f $ **FLOATING
C16 a_n440_n514# VSS 0.59507f $ **FLOATING
C17 a_n440_286# VSS 0.59511f $ **FLOATING
C18 a_n441_1087# VSS 0.59126f $ **FLOATING
C19 a_n441_1887# VSS 0.60422f $ **FLOATING
C20 a_n441_2690# VSS 0.58987f $ **FLOATING
.ends

