* NGSPICE file created from LELO_EX.ext - technology: sky130A

.subckt JNWATR_NCH_4C5F0 D G S B a_160_778# a_160_n22# a_1056_n40#
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X1 S G D B sky130_fd_pr__nfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
.ends

.subckt LELO_EX IBPS_5U IBNS_20U VSS
XJNWATR_NCH_4C5F0_0 IBNS_20U IBPS_5U VSS VSS JNWATR_NCH_4C5F0_1/a_160_n22# JNWATR_NCH_4C5F0_0/a_160_n22#
+ JNWATR_NCH_4C5F0_0/a_1056_n40# JNWATR_NCH_4C5F0
XJNWATR_NCH_4C5F0_1 IBNS_20U IBPS_5U VSS VSS JNWATR_NCH_4C5F0_2/a_160_n22# JNWATR_NCH_4C5F0_1/a_160_n22#
+ JNWATR_NCH_4C5F0_1/a_1056_n40# JNWATR_NCH_4C5F0
XJNWATR_NCH_4C5F0_2 IBPS_5U IBPS_5U VSS VSS JNWATR_NCH_4C5F0_3/a_160_n22# JNWATR_NCH_4C5F0_2/a_160_n22#
+ VSS JNWATR_NCH_4C5F0
XJNWATR_NCH_4C5F0_3 IBNS_20U IBPS_5U VSS VSS JNWATR_NCH_4C5F0_4/a_160_n22# JNWATR_NCH_4C5F0_3/a_160_n22#
+ VSS JNWATR_NCH_4C5F0
XJNWATR_NCH_4C5F0_4 IBNS_20U IBPS_5U VSS VSS JNWATR_NCH_4C5F0_4/a_160_778# JNWATR_NCH_4C5F0_4/a_160_n22#
+ VSS JNWATR_NCH_4C5F0
.ends

