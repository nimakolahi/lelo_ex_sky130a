** sch_path: /home/n.mahmoudi/pro/aicex/ip/lelo_ex_sky130a/design/LELO_EX_SKY130A/LELO_EX.sch
.subckt LELO_EX IBPS_5U VSS IBNS_20U
*.ipin IBPS_5U
*.ipin VSS
*.opin IBNS_20U
xo<3> IBNS_20U IBPS_5U VSS VSS JNWATR_NCH_4C5F0
xo<2> IBNS_20U IBPS_5U VSS VSS JNWATR_NCH_4C5F0
xo<1> IBNS_20U IBPS_5U VSS VSS JNWATR_NCH_4C5F0
xo<0> IBNS_20U IBPS_5U VSS VSS JNWATR_NCH_4C5F0
xi IBPS_5U IBPS_5U VSS VSS JNWATR_NCH_4C5F0
.ends

* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym # of pins=4
** sym_path: /home/n.mahmoudi/pro/aicex/ip/lelo_ex_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym
** sch_path: /home/n.mahmoudi/pro/aicex/ip/lelo_ex_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sch
.subckt JNWATR_NCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
